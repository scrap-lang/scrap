module main

struct File {
mut:
	stmts []Stmt
}

fn parse(input string) ?File {
	// TODO: this.
}

fn main() {
	code = "let foo = 10"
}
